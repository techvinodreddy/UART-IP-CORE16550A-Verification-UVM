package test_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"
  
  `include "xtn.sv"
  `include "agt_config.sv"
  `include "env_config.sv"

  `include "seqs.sv"
  `include "seqr.sv"
  `include "drv.sv"
  `include "mon.sv"
  `include "agt.sv"
  `include "agt_top.sv"

  `include "v_seqr.sv"
  `include "v_seqs.sv"
  `include "scoreboard.sv"

  `include "env.sv"
  `include "test.sv"
endpackage
