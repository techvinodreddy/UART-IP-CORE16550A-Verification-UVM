`define DBS 8  // Data Bus Modes data_in, data_out size 8 or 32
`define ADDR 5 // Address register size 3 or 5
`define SEL 4  // Select Signal
